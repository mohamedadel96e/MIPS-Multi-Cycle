LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
ENTITY MUX_3to1 IS
  GENERIC (N : INTEGER := 32);
  PORT (
    Sel : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    In0 : IN STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
    In1 : IN STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
    In2 : IN STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
    OutMux : OUT STD_LOGIC_VECTOR(N - 1 DOWNTO 0)
  );
END ENTITY;

ARCHITECTURE Behavioral OF MUX_3to1 IS
BEGIN
  OutMux <= In0 WHEN Sel = "00" ELSE
    In1 WHEN Sel = "01" ELSE
    In2;
END Behavioral;