library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity MultiCycleMips is 
  port (
    clk : in std_logic;
    reset : in std_logic
  );
end entity;